CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 110 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 76 128 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89884e-315 0
0
2 +V
167 200 247 0 1 3
0 2
0
0 0 54256 180
2 5V
10 -2 24 6
3 V10
6 -12 27 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
391 0 0
2
43530.4 0
0
2 +V
167 321 248 0 1 3
0 3
0
0 0 54256 180
2 5V
7 -2 21 6
2 V9
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3124 0 0
2
43530.4 0
0
2 +V
167 474 244 0 1 3
0 4
0
0 0 54256 180
2 5V
7 -2 21 6
2 V8
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3421 0 0
2
43530.4 0
0
6 74112~
219 474 219 0 7 32
0 5 22 23 22 4 25 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
8157 0 0
2
43530.4 0
0
2 +V
167 716 252 0 1 3
0 6
0
0 0 54256 180
2 5V
7 -2 21 6
2 V7
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5572 0 0
2
43530.4 0
0
2 +V
167 721 234 0 1 3
0 2
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
43530.4 0
0
2 +V
167 716 161 0 1 3
0 7
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
43530.4 0
0
2 +V
167 474 150 0 1 3
0 5
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
43530.4 0
0
2 +V
167 321 153 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
43530.4 0
0
9 CC 7-Seg~
183 1163 139 0 18 19
10 20 19 18 17 16 15 14 26 27
1 0 0 1 0 1 1 2 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3472 0 0
2
5.89884e-315 5.26354e-315
0
2 +V
167 200 139 0 1 3
0 13
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.89884e-315 5.30499e-315
0
6 74LS48
188 807 303 0 14 29
0 12 11 10 9 28 29 14 15 16
17 18 19 20 30
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.89884e-315 5.32571e-315
0
9 2-In AND~
219 548 52 0 3 22
0 22 11 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4597 0 0
2
5.89884e-315 5.34643e-315
0
9 2-In AND~
219 380 44 0 3 22
0 9 10 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3835 0 0
2
5.89884e-315 5.3568e-315
0
7 Pulser~
4 82 261 0 10 12
0 31 32 23 33 0 0 5 5 4
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3670 0 0
2
5.89884e-315 5.36716e-315
0
6 74112~
219 716 230 0 7 32
0 7 21 23 21 6 34 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
5616 0 0
2
5.89884e-315 5.37752e-315
0
6 74112~
219 321 224 0 7 32
0 8 9 23 9 3 35 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
9323 0 0
2
5.89884e-315 5.39306e-315
0
6 74112~
219 200 224 0 7 32
0 13 24 23 24 2 36 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
317 0 0
2
5.89884e-315 5.39824e-315
0
35
1 5 2 0 0 4224 0 2 19 0 0 2
200 232
200 236
1 5 3 0 0 4224 0 3 18 0 0 2
321 233
321 236
1 5 4 0 0 4224 0 4 5 0 0 2
474 229
474 231
1 1 5 0 0 4224 0 5 9 0 0 2
474 156
474 159
1 5 6 0 0 4224 0 6 17 0 0 2
716 237
716 242
1 1 7 0 0 4224 0 8 17 0 0 2
716 170
716 167
1 1 8 0 0 4224 0 10 18 0 0 2
321 162
321 161
4 0 9 0 0 12416 0 13 0 0 29 5
775 294
767 294
767 359
237 359
237 188
0 3 10 0 0 12416 0 0 13 26 0 6
349 174
407 174
407 347
756 347
756 285
775 285
0 2 11 0 0 8320 0 0 13 22 0 6
511 179
590 179
590 335
745 335
745 276
775 276
7 1 12 0 0 8320 0 17 13 0 0 4
740 194
766 194
766 267
775 267
1 1 13 0 0 4224 0 12 19 0 0 2
200 148
200 161
7 7 14 0 0 8320 0 11 13 0 0 3
1178 175
1178 267
839 267
8 6 15 0 0 4224 0 13 11 0 0 3
839 276
1172 276
1172 175
9 5 16 0 0 4224 0 13 11 0 0 3
839 285
1166 285
1166 175
10 4 17 0 0 4224 0 13 11 0 0 3
839 294
1160 294
1160 175
11 3 18 0 0 4224 0 13 11 0 0 3
839 303
1154 303
1154 175
12 2 19 0 0 4224 0 13 11 0 0 3
839 312
1148 312
1148 175
13 1 20 0 0 4224 0 13 11 0 0 3
839 321
1142 321
1142 175
4 0 21 0 0 4096 0 17 0 0 21 3
692 212
611 212
611 186
3 2 21 0 0 8320 0 14 17 0 0 4
569 52
611 52
611 194
692 194
2 7 11 0 0 16 0 14 5 0 0 4
524 61
511 61
511 183
498 183
1 0 22 0 0 4096 0 14 0 0 25 3
524 43
412 43
412 96
0 4 22 0 0 0 0 0 5 25 0 4
412 187
413 187
413 201
450 201
3 2 22 0 0 8320 0 15 5 0 0 6
401 44
412 44
412 187
412 187
412 183
450 183
2 7 10 0 0 0 0 15 18 0 0 4
356 53
349 53
349 188
345 188
1 0 9 0 0 0 0 15 0 0 28 3
356 35
282 35
282 188
4 0 9 0 0 0 0 18 0 0 29 3
297 206
282 206
282 188
7 2 9 0 0 0 0 19 18 0 0 2
224 188
297 188
3 0 23 0 0 12416 0 17 0 0 31 4
686 203
672 203
672 252
418 252
3 0 23 0 0 0 0 5 0 0 32 6
444 192
444 227
418 227
418 252
291 252
291 251
3 0 23 0 0 0 0 18 0 0 35 3
291 197
291 251
121 251
1 0 24 0 0 8320 0 1 0 0 34 3
88 128
138 128
138 188
2 4 24 0 0 0 0 19 19 0 0 4
176 188
137 188
137 206
176 206
3 3 23 0 0 0 0 19 16 0 0 5
170 197
170 251
121 251
121 252
106 252
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
